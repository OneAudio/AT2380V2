OSC_inst : OSC PORT MAP (
		oscena	 => oscena_sig,
		osc	 => osc_sig
	);
